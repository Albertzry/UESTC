module INSTMEM(Addr,Inst);
input[31:0]Addr;
output[31:0]Inst;
wire[31:0]Rom[31:0];
assign Rom[5'h00]=32'b001000_00000_00001_0000_0000_0000_0110;//addi $1,$0,6 $1=6
assign Rom[5'h01]=32'b001101_00000_00010_0000_0000_0000_1100;//ori $2,$0,12 $2=12
assign Rom[5'h02]=32'b001100_00001_00011_1111_1111_1111_1111;//andi $3,$1,65535 $3=6
assign Rom[5'h03]=32'b001110_00010_00100_0000_0000_0000_1111;//xori $4,$2,15 $4=3
assign Rom[5'h04]=32'hXXXXXXXX;
assign Rom[5'h05]=32'b000000_00001_00010_00101_00000_100000;//and $5,$1,$2 $5=18
assign Rom[5'h06]=32'b000000_00010_00001_00110_00000_100010;//sub $6,$2,$1 $6=6
assign Rom[5'h07]=32'b000000_00001_00010_00111_00000_100100;//and $7,$1,$2 $7=4
assign Rom[5'h08]=32'b000000_00001_00100_01000_00000_100101;//or $8,$1,$4 $8=7
assign Rom[5'h09]=32'b000000_00001_00010_01001_00000_100110;//xor $9,$1,$2 $9=10
assign Rom[5'h0A]=32'b000000_00000_00001_01010_00010_000000;//sll $10,$1 2 $10=24
assign Rom[5'h0B]=32'b000000_00000_00010_01011_00010_000010;//srl $11,$2 2 $11=3
assign Rom[5'h0C]=32'b000000_00000_00001_01100_00001_000011;//sra $12,$1 1 $12=3
assign Rom[5'h0D]=32'hXXXXXXXX;
assign Rom[5'h0E]=32'b101011_01000_00010_0000000000001010;//sw $1 10($8) memory[$8+10]=6
assign Rom[5'h0F]=32'b100011_01000_01101_0000000000001010;//lw $13 10($8) $13=12
assign Rom[5'h10]=32'b000100_00001_00011_0000000000000010;//beq $1 $3 2
assign Rom[5'h11]=32'hXXXXXXXX;
assign Rom[5'h12]=32'hXXXXXXXX;
assign Rom[5'h13]=32'b000000_01001_01000_01110_00000_100000;//and $14 $9 $8 $14=17
assign Rom[5'h14]=32'b000101_00001_00010_0000000000000011;//	bne $1 $2 3
assign Rom[5'h15]=32'hXXXXXXXX;
assign Rom[5'h16]=32'hXXXXXXXX;
assign Rom[5'h17]=32'hXXXXXXXX;
assign Rom[5'h18]=32'b001111_00000_01111_0000000000000000;//lui $15 
assign Rom[5'h19]=32'b000011_00000000000000000000011100;//jal
assign Rom[5'h1A]=32'b000010_00000000000000000000011100;//j
assign Rom[5'h1B]=32'hXXXXXXXX;
assign Rom[5'h1C]=32'b000000_00000_00000_00000_00000_001000;//jr $0
assign Rom[5'h1D]=32'hXXXXXXXX;		
assign Rom[5'h1E]=32'hXXXXXXXX;
assign Rom[5'h1F]=32'hXXXXXXXX;
assign Inst=Rom[Addr[6:2]];
endmodule
